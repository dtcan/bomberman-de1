module bomberman_control
endmodule
