module bomberman();
endmodule
