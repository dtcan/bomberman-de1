module bomberman_datapath
endmodule
